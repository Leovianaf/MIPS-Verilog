// Universidade Federal Rural de Pernambuco
// 2023.1
// Arquitetura e Organização de Computadores - 2ªVA
// Alunos:
// Beatriz Pereira, Leonardo Viana, Paloma Raissa, Ricardo Zaidan
// -----------------------------

module pc(nextPC, pc, clock);

	// Declaração de entradas e saída
	input clock;
	input wire [31:0] nextPC;
	output reg [31:0] pc;
	
	// Declaração de flag
	reg reset;

	// Inicializando reset = 0 e pc = 0
	initial begin
		reset = 0;
		pc = 32'b0;
	end

	// Atribuição síncrona. Se reset == 1, pc recebe o valor de nextPC. Se reset == 0, PC é zerado
	always @(posedge clock) begin
		if(reset) begin
			pc = nextPC;
		end else begin
			pc = 32'b0;
			reset = 1;
		end
	end
endmodule
